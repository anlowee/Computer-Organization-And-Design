`timescale 1ns/1ps
module alu_test;
    reg[31:0] a, b;
    reg[2:0] opcode;
    wire[2:0] d;
    wire[31:0] c;

    parameter sla = 3'b000,
        sra = 3'b001,
        add = 3'b010,
        sub = 3'b011,
        mul = 3'b100,
        andd = 3'b101,
        ord = 3'b110,
        notd = 3'b111;
    
    alu testalu(a, b, opcode, c, d);

    initial
    begin
        #10 a = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            b = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            opcode = mul;
        #10 a = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            b = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            opcode = mul;
        #10 a = 32'b1111_1111_1111_1110_0000_0000_0000_0000;
            b = 32'b1111_1111_1111_1110_0000_0000_0000_0000;
            opcode = mul;
        #10 a = 32'b1111_1111_1111_1111_1111_1111_1111_1110;
            b = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            opcode = mul;
        #10 a = 32'b1111_1111_1111_1110_0000_0000_0000_0000;
            b = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            opcode = mul;

        #10 $finish;
    end


endmodule
